module Execute (
    
);
    
endmodule